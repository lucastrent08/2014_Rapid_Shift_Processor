----------------------------------------------------------------------------------
-- Company: Bryant Electric Motors/University of Massachusetts Dartmouth
-- Department: Electrical and Computer Engineering
-- Engineer: Lucas Trent
-- Create Date:    March 2014
-- Module Name:    FPU
-- Project Name: 	 CISC 04
-- Target Devices: Spartan-3E
-- Tool versions:	 Xilinx ISE 9.2-- Description: CCU Microprogram ROM.
---------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity microprogram_rom is
   port(
      clk: in std_logic;
      address : in std_logic_vector (7 downto 0);
		output : out std_logic_vector (69 downto 0)
   );
end microprogram_rom;

architecture Behavioral of microprogram_rom is
	
	signal output_reg : std_logic_vector (69 downto 0) := (OTHERS => '0');
   type rom_type is array (0 to 2**8-1)
        of std_logic_vector (69 downto 0);
   signal rom: rom_type := (
--CCR: BRA          LC   MASK              BS  AS PCU: CI  INSTR   OE SSCU: CEM CI   SHIFT  INSTR    S   Ceu ALU: Dest   Fctn   Src   IDB MEM: VMA RW  DBB IR
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00001"&'0'&     '1'&"00"&"0000"&"000000"&'0'&'1'&     "0000"&"0000"&"000"&"000"&   '1'&'1'&'1'&'1', -- $00
		"00000000001"&'0'&"0000000000000000"&'0'&'0' &   '1'&"00001"&'0'&     '1'&"00"&"0000"&"000000"&'0'&'0'&     "0000"&"0000"&"000"&"000"&   '1'&'1'&'1'&'0', -- $01
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $02
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $03
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"10100"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "0000"&"0000"&"000"&"110"&   '0'&'1'&'1'&'1', -- $04
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $05
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $06
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $07
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '1'&"10100"&'0'&     '1'&"00"&"0000"&"000000"&'0'&'1'&     "1100"&"0110"&"000"&"110"&   '0'&'1'&'0'&'1', -- $08
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $09
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'1'&     '0'&"01"&"0000"&"000110"&'1'&'1'&     "1111"&"0001"&"000"&"101"&   '0'&'1'&'1'&'1', -- $0A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $0B
		"00000000000"&'0'&"0000000000001111"&'0'&'0' &   '0'&"01111"&'1'&     '0'&"01"&"1010"&"000110"&'1'&'1'&     "1111"&"0001"&"100"&"101"&   '0'&'1'&'1'&'1', -- $0C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $0D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $0E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $0F
		"00000000000"&'0'&"0000000000001111"&'0'&'0' &   '0'&"11111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0110"&"100"&"101"&   '0'&'1'&'1'&'1', -- $10
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $11
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $12
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $13
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"11111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0110"&"100"&"000"&   '0'&'1'&'0'&'1', -- $14
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $15
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $16
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $17
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"11111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0110"&"000"&"001"&   '0'&'1'&'1'&'1', -- $18
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"11111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'0'&'0'&'1', -- $19
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $1A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $1B
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $1C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $1D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $1E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $1F
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '1'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "0000"&"0000"&"000"&"000"&   '0'&'1'&'0'&'1', -- $20
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00001"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0011"&"000"&"001"&   '1'&'0'&'1'&'1', -- $21
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $22
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $23
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $24
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $25
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $26
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $27
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01100"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0110"&"000"&"001"&   '0'&'1'&'1'&'1', -- $28
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $29
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $2A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $2B
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $2C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $2D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $2E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $2F
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01101"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0110"&"100"&"010"&   '0'&'1'&'1'&'1', -- $30
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $31
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $32
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $33
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $34
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $35
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $36
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $37
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'1'&'1'&'1', -- $38
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "0110"&"0011"&"100"&"000"&   '0'&'1'&'0'&'1', -- $39
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0110"&"000"&"000"&   '0'&'1'&'1'&'1', -- $3A
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"010"&"000"&   '1'&'0'&'0'&'1', -- $3B
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $3C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $3D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $3E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $3F
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '1'&"01010"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '0'&'1'&'0'&'1', -- $40
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00010"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'1'&'1'&'1', -- $41
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'1'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1111"&"0011"&"100"&"001"&   '0'&'1'&'1'&'1', -- $42
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $43
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $44
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $45
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $46
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $47
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $48
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $49
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $4A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $4B
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $4C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $4D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $4E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $4F
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0110"&"000"&"001"&   '0'&'1'&'1'&'1', -- $50
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $51
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $52
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $53
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0011"&"000"&"001"&   '0'&'1'&'1'&'1', -- $54
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0011"&"000"&"001"&   '0'&'1'&'1'&'1', -- $55
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $56
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $57
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $58
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $59
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $5A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $5B
		"00000000111"&'0'&"0000000000001111"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"101"&   '0'&'1'&'1'&'1', -- $5C
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'0'&'0'&'1', -- $5D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $5E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $5F
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $60
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $61
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $62
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $63
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $64
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $65
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $66
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $67
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '1'&"00001"&'1'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1111"&"1100"&"100"&"000"&   '0'&'1'&'0'&'1', -- $68
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $69
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $6A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $6B
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0110"&"000"&"001"&   '1'&'1'&'1'&'1', -- $6C
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "0110"&"0110"&"100"&"000"&   '0'&'1'&'0'&'1', -- $6D
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'1'&'1'&'1', -- $6E
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'1'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1111"&"0001"&"100"&"001"&   '0'&'1'&'1'&'1', -- $6F
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '1'&"00010"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"000"&   '0'&'1'&'0'&'1', -- $70
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00010"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'1'&'1'&'1', -- $71
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'1'&     '0'&"00"&"0000"&"000110"&'1'&'1'&     "0110"&"0011"&"100"&"000"&   '0'&'1'&'0'&'1', -- $72
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"010"&"001"&   '0'&'1'&'1'&'1', -- $73
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00010"&'0'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'0'&'0'&'1', -- $74
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $75
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $76
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $77
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $78
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $79
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $7A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $7B
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $7C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $7D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $7E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $7F
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0110"&"000"&"001"&   '1'&'1'&'1'&'1', -- $80
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "0110"&"0110"&"100"&"000"&   '0'&'1'&'0'&'1', -- $81
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'1'&'1'&'1', -- $82
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'1'&     '0'&"00"&"0000"&"000110"&'1'&'1'&     "0110"&"0011"&"110"&"000"&   '0'&'1'&'0'&'1', -- $83
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"010"&"001"&   '0'&'1'&'1'&'1', -- $84
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1100"&"0100"&"000"&"001"&   '1'&'0'&'0'&'1', -- $85
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $86
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $87
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $88
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $89
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $8A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $8B
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00011"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0110"&"000"&"001"&   '1'&'1'&'1'&'1', -- $8C
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01100"&'0'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1100"&"0100"&"000"&"000"&   '0'&'1'&'0'&'1', -- $8D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $8E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $8F
		"00000000110"&'0'&"0000000000001111"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "1100"&"0100"&"000"&"101"&   '0'&'1'&'1'&'1', -- $90
		"00000000100"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'1'&     '0'&"00"&"0000"&"000110"&'1'&'0'&     "0000"&"0100"&"000"&"001"&   '0'&'1'&'1'&'1', -- $91
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"001"&   '0'&'1'&'1'&'1', -- $92
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $93
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $94
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $95
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $96
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $97
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $98
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $99
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $9A
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $9B
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $9C
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $9D
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $9E
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $9F
		"00000000001"&'1'&"0000000000000000"&'0'&'0' &   '1'&"00001"&'0'&     '1'&"00"&"0000"&"000101"&'1'&'0'&     "1111"&"0001"&"100"&"111"&   '0'&'1'&'0'&'1', -- $A0
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"10100"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"000"&   '0'&'1'&'1'&'1', -- $A1
		
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '1'&"00001"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"000"&   '1'&'1'&'0'&'1', -- $A2
		"00000000111"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01010"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0100"&"000"&"000"&   '0'&'1'&'0'&'1', -- $A3
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"00010"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1111"&"0100"&"000"&"001"&   '1'&'0'&'0'&'1', -- $A4
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $A5	
		
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"10001"&'0'&     '0'&"00"&"0000"&"000000"&'0'&'0'&     "1100"&"0100"&"000"&"000"&   '1'&'1'&'0'&'1', -- $A6
		
		"00000000000"&'0'&"0000000000000000"&'0'&'0' &   '0'&"01111"&'0'&     '0'&"01"&"0000"&"000000"&'0'&'0'&     "1111"&"0100"&"000"&"000"&   '0'&'1'&'1'&'1', -- $A7
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $A8
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $A9
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $AA
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $AB
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $AC
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $AD
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $AE
		"0000000000000000000000000000000000000000000000000000000000000000000000", -- $AF
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000000000"
		);
begin
	-- read cycle
   process(clk)
   begin
     if (clk'event and clk = '1') then
        output_reg <= rom(to_integer(unsigned(address)));
     end if;
   end process;
	output <= output_reg;

end Behavioral;
